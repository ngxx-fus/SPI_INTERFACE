`include "sender_receiver.v"
`include "control.v"
`include "status.v"

module SPI(
	input MS_MODE,
	input CLK,
	input CLR,
	input READ,
	input WRITE,
	input  [7:0] CONTROL,
	output [7:0] STATUS,
	input  [7:0] INCOMING_DATA,
	output [7:0] OUTCOMING_DATA,
	input MISO,
	output MOSI,
	inout CS,
	inout S_CLK
);
	wire HIGH, LOW;

	wire LOCAL_CLK;
	wire SENDER_CLK;
	wire SENDER_CLR;
	wire SENDER_WRITE;
	wire TE;
	wire SENDER_REG_FULL;
	wire SENDER_EMPTY_STATE;
	
	wire RECEIVER_CLK;
	wire RECEIVER_CLR;
	wire RECEIVER_READ;
	wire RE;
	wire RECEIVER_FULL_STATE;
	wire RECEIVER_EMPTY_STATE;

	wire [7:0] SENDER_BUFFER_DATA_I;
	wire [7:0] SENDER_BUFFER_DATA_O;
	wire       SENDER_BUFFER_SH_LD;

	wire [7:0] RECEIVER_BUFFER_DATA_I;
	wire [7:0] RECEIVER_BUFFER_DATA_O;
	wire       RECEIVER_BUFFER_SH_LD;

	wire CONNECTION_FAILED_STATE;
	wire CS_CONTROL;
	wire LOCAL_MOSI;

	//since the 8bit register is PIPO,
	//so it can only FULL or EMPTY :v
	wire SENDER_BUFFER_FULL_STATE;
	SHIFT_REGISTER_8BIT SENDER_BUFFER(
		.CLK(LOW),
		.CLR(CLR),
		.P_DATA_IN(SENDER_BUFFER_DATA_I),
		.SH_LD(SENDER_BUFFER_SH_LD),
		.P_DATA_OUT(SENDER_BUFFER_DATA_O)
	);

	wire RECEIVER_BUFFER_FULL_STATE;	
	SHIFT_REGISTER_8BIT RECEIVER_BUFFER(
		.CLK(LOW),
		.CLR(CLR),
		.P_DATA_IN(RECEIVER_BUFFER_DATA_I),
		.SH_LD(RECEIVER_BUFFER_SH_LD),
		.P_DATA_OUT(RECEIVER_BUFFER_DATA_O)
	);
	
	SENDER sender(
		.CLK(SENDER_CLK),
		.CLR(SENDER_CLR),
		.WRITE(SENDER_WRITE),
		.TE(TE),
		.FULL_STATE(SENDER_FULL_STATE),
		.EMPTY_STATE(SENDER_EMPTY_STATE),
		.DATA(SENDER_BUFFER_DATA_O),
		.MOSI(LOCAL_MOSI)
	);
	RECEIVER receiver(
		.CLK(RECEIVER_CLK),
		.CLR(RECEIVER_CLR),
		.READ(RECEIVER_READ),
		.RE(RE),
		.FULL_STATE(RECEIVER_FULL_STATE),
		.EMPTY_STATE(RECEIVER_EMPTY_STATE),
		.DATA(RECEIVER_BUFFER_DATA_I),
		.MISO(MISO)
	);
	STATUS_COMBINATION status(
		//command signal
		.S_CLK(S_CLK),
		.CLR(CLR),
		.SENDER_WRITE(SENDER_WRITE),
		//buffer
		.SENDER_BUFFER_SH_LD(SENDER_BUFFER_SH_LD),
		.SENDER_BUFFER_FULL_STATE(SENDER_BUFFER_FULL_STATE),
		.RECEIVER_BUFFER_SH_LD(RECEIVER_BUFFER_SH_LD),
		.RECEIVER_BUFFER_FULL_STATE(RECEIVER_BUFFER_FULL_STATE),
		//status of sender
		.SENDER_FULL_STATE(SENDER_FULL_STATE),
		.SENDER_EMPTY_STATE(SENDER_EMPTY_STATE),
		//status of receiver
		.RECEIVER_FULL_STATE(RECEIVER_FULL_STATE),
		.RECEIVER_EMPTY_STATE(RECEIVER_EMPTY_STATE),
		.STATUS(STATUS),
		.CONNECTION_FAILED_STATE(CONNECTION_FAILED_STATE)
	);
	
	CONTROL_COMBINATION control(
		.MS_MODE(MS_MODE),
		.CLK(LOCAL_CLK),
		.CLR(CLR),
		.CONTROL(CONTROL),
		.WRITE(WRITE),
		.READ(READ),
		.SENDER_BUFFER_FULL_STATE(SENDER_BUFFER_FULL_STATE),
		.SENDER_BUFFER_SH_LD(SENDER_BUFFER_SH_LD),
		.RECEIVER_BUFFER_FULL_STATE(RECEIVER_BUFFER_FULL_STATE),
		.RECEIVER_BUFFER_SH_LD(RECEIVER_BUFFER_SH_LD),
		.SENDER_CLK(SENDER_CLK),
		.SENDER_CLR(SENDER_CLR),
		.SENDER_FULL_STATE(SENDER_FULL_STATE),
		.SENDER_EMPTY_STATE(SENDER_EMPTY_STATE),
		.SENDER_WRITE(SENDER_WRITE),
		.TE(TE),
		.RECEIVER_CLK(RECEIVER_CLK),
		.RECEIVER_CLR(RECEIVER_CLR),
		.RECEIVER_FULL_STATE(RECEIVER_FULL_STATE),
		.RECEIVER_EMPTY_STATE(RECEIVER_EMPTY_STATE),
		.RE(RE),
		.RECEIVER_READ(RECEIVER_READ),
		.CS(CS_CONTROL)
	);

	assign MOSI = (MS_MODE==HIGH)?(LOCAL_MOSI):((CS==HIGH)?1'bz:LOCAL_MOSI);
	assign LOCAL_CLK = (MS_MODE==HIGH)?(CLK):(S_CLK);
	assign S_CLK = (MS_MODE == HIGH)?(CLK & (~CS)):(1'bz);
	assign OUTCOMING_DATA = (READ==HIGH)?RECEIVER_BUFFER_DATA_O:8'hzz;
	assign SENDER_BUFFER_DATA_I = INCOMING_DATA;
	assign CONNECTION_FAILED_STATE = ((CS != 1 && CS!=0) 
	                                ||(MISO != 1 && MISO!=0) 
	                                ||(S_CLK != 1 && S_CLK!=0)  )?HIGH:LOW;
	assign CS = (MS_MODE==HIGH)?(CS_CONTROL):1'bz;
	assign LOW = 1'b0;
	assign HIGH = 1'b1;
endmodule
